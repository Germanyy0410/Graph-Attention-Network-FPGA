module softmax #(

)(

);
endmodule