`define SIMULATION            1

// `define CORA                  1
// `define CITESEER              1
// `define PUBMED                1

// `define VIVADO                1

// `define PASSED                1
`define FAILED                1