// ==================================================================
// File name  : gat_define.sv
// Project    : Graph Attention Network Accelerator on FPGA
// Function   :
// -- All defines used in the project
// -- Used to switch between Simulation, Synthesis, Dataset, etc.
// Author     : @Germanyy0410
// ==================================================================

// `define SIMULATION            1

// `define CORA                  1
// `define CITESEER              1
// `define PUBMED                1

// `define VIVADO                1

// `define PASSED                1
`define FAILED                1