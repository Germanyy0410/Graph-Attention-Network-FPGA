module top #(

)(

);
endmodule