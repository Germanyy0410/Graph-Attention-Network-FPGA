module SPV #(

)(

);
endmodule