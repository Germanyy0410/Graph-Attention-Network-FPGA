module SPMM #(

)(

);
endmodule