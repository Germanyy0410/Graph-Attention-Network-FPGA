package define_pkg;
  `define SIMULATION            1

  // `define CORA_DATASET_EN       1
  // `define CITESEER_DATASET_EN   1
  // `define PUBMED_DATASET_EN     1
endpackage