module DMVM #(

)(

);
endmodule