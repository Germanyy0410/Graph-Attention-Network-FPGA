module SP_PE #(
  //* ====================== parameter ========================
  parameter DATA_WIDTH            = 8,
  parameter WH_DATA_WIDTH         = 12,
  parameter DMVM_DATA_WIDTH       = 19,
  parameter SM_DATA_WIDTH         = 108,
  parameter SM_SUM_DATA_WIDTH     = 108,
  parameter ALPHA_DATA_WIDTH      = 32,
  parameter NEW_FEATURE_WIDTH     = 32,

  parameter H_NUM_SPARSE_DATA     = 242101,
  parameter TOTAL_NODES           = 13264,
  parameter NUM_FEATURE_IN        = 1433,
  parameter NUM_FEATURE_OUT       = 16,
  parameter NUM_SUBGRAPHS         = 2708,
  parameter MAX_NODES             = 168,

  parameter COEF_DEPTH            = 500,
  parameter ALPHA_DEPTH           = 500,
  parameter DIVIDEND_DEPTH        = 500,
  parameter DIVISOR_DEPTH         = 500,
  //* =========================================================

  //* ====================== localparams ======================
  // -- [BRAM]
  localparam H_DATA_DEPTH         = H_NUM_SPARSE_DATA,
  localparam NODE_INFO_DEPTH      = TOTAL_NODES,
  localparam WEIGHT_DEPTH         = NUM_FEATURE_OUT * NUM_FEATURE_IN + NUM_FEATURE_OUT * 2,
  localparam WH_DEPTH             = TOTAL_NODES,
  localparam A_DEPTH              = NUM_FEATURE_OUT * 2,
  localparam NUM_NODES_DEPTH      = NUM_SUBGRAPHS,
  localparam NEW_FEATURE_DEPTH    = NUM_SUBGRAPHS * NUM_FEATURE_OUT,

  // -- [H]
  localparam H_NUM_OF_ROWS        = TOTAL_NODES,
  localparam H_NUM_OF_COLS        = NUM_FEATURE_IN,

  // -- [H] data
  localparam COL_IDX_WIDTH        = $clog2(H_NUM_OF_COLS),
  localparam H_DATA_WIDTH         = DATA_WIDTH + COL_IDX_WIDTH,
  localparam H_DATA_ADDR_W        = $clog2(H_DATA_DEPTH),

  // -- [H] node_info
  localparam ROW_LEN_WIDTH        = $clog2(H_NUM_OF_COLS),
  localparam NUM_NODE_WIDTH       = $clog2(MAX_NODES),
  localparam FLAG_WIDTH           = 1,
  localparam NODE_INFO_WIDTH      = ROW_LEN_WIDTH + NUM_NODE_WIDTH + FLAG_WIDTH,
  localparam NODE_INFO_ADDR_W     = $clog2(NODE_INFO_DEPTH),

  // -- [W]
  localparam W_NUM_OF_ROWS        = NUM_FEATURE_IN,
  localparam W_NUM_OF_COLS        = NUM_FEATURE_OUT,
  localparam W_ROW_WIDTH          = $clog2(W_NUM_OF_ROWS),
  localparam W_COL_WIDTH          = $clog2(W_NUM_OF_COLS),
  localparam WEIGHT_ADDR_W        = $clog2(WEIGHT_DEPTH),
  localparam MULT_WEIGHT_ADDR_W   = $clog2(W_NUM_OF_ROWS),

  // -- [WH]
  localparam DOT_PRODUCT_SIZE     = H_NUM_OF_COLS,
  localparam WH_ADDR_W            = $clog2(WH_DEPTH),
  localparam WH_RESULT_WIDTH      = WH_DATA_WIDTH * W_NUM_OF_COLS,
  localparam WH_WIDTH             = WH_DATA_WIDTH * W_NUM_OF_COLS + NUM_NODE_WIDTH + FLAG_WIDTH,

  // -- [A]
  localparam A_ADDR_W             = $clog2(A_DEPTH),
  localparam HALF_A_SIZE          = A_DEPTH / 2,
  localparam A_INDEX_WIDTH        = $clog2(A_DEPTH),

  // -- [DMVM]
  localparam DMVM_PRODUCT_WIDTH   = $clog2(HALF_A_SIZE),
  localparam COEF_W               = DATA_WIDTH * MAX_NODES,
  localparam ALPHA_W              = ALPHA_DATA_WIDTH * MAX_NODES,
  localparam NUM_NODE_ADDR_W      = $clog2(NUM_NODES_DEPTH),
  localparam NUM_STAGES           = $clog2(NUM_FEATURE_OUT) + 1,
  localparam COEF_DELAY_LENGTH    = NUM_STAGES + 1,

  // -- [SOFTMAX]
  localparam SOFTMAX_WIDTH        = MAX_NODES * DATA_WIDTH + NUM_NODE_WIDTH,
  localparam SOFTMAX_DEPTH        = NUM_SUBGRAPHS,
  localparam SOFTMAX_ADDR_W       = $clog2(SOFTMAX_DEPTH),
  localparam WOI                  = 1,
  localparam WOF                  = ALPHA_DATA_WIDTH - WOI,
  localparam DL_DATA_WIDTH        = $clog2(WOI + WOF + 3) + 1,
  localparam DIVISOR_FF_WIDTH     = NUM_NODE_WIDTH + SM_SUM_DATA_WIDTH,

  // -- [AGGREGATOR]
  localparam AGGR_WIDTH           = MAX_NODES * ALPHA_DATA_WIDTH + NUM_NODE_WIDTH,
  localparam AGGR_DEPTH           = NUM_SUBGRAPHS,
  localparam AGGR_ADDR_W          = $clog2(AGGR_DEPTH),
  localparam AGGR_MULT_W          = WH_DATA_WIDTH + 32,

  // -- [NEW FEATURE]
  localparam NEW_FEATURE_ADDR_W   = $clog2(NEW_FEATURE_DEPTH)
  //* =========================================================
)(
  input                             clk                     ,
  input                             rst_n                   ,

  input                             spmm_vld_i              ,
  input                             pe_vld_i                ,
  output                            pe_rdy_o                ,

  input   [COL_IDX_WIDTH-1:0]       col_idx_i               ,
  input   [DATA_WIDTH-1:0]          val_i                   ,

  input   [ROW_LEN_WIDTH-1:0]       row_len_i               ,
  input   [NUM_NODE_WIDTH-1:0]      num_node_i              ,
  input                             src_flag_i              ,

  output  [NUM_NODE_WIDTH-1:0]      num_node_o              ,
  output                            src_flag_o              ,

  input   [DATA_WIDTH-1:0]          wgt_dout                ,
  output  [MULT_WEIGHT_ADDR_W-1:0]  wgt_addrb               ,

  output  [ROW_LEN_WIDTH:0]         cnt_reg                 ,

  output  [WH_DATA_WIDTH-1:0]       res_o
);

  //* =================== logic declaration ===================
  logic                               spmm_vld_q1         ;

  logic         [COL_IDX_WIDTH-1:0]   col_idx_reg         ;
  logic         [DATA_WIDTH-1:0]      val_reg             ;
  logic         [ROW_LEN_WIDTH-1:0]   row_len_reg         ;
  // -- [pe_rdy] logic
  logic                               pe_rdy              ;
  logic                               pe_rdy_reg          ;
  // -- [res] logic
  logic signed  [WH_DATA_WIDTH-1:0]   res                 ;
  logic signed  [WH_DATA_WIDTH-1:0]   res_reg             ;

  logic signed  [WH_DATA_WIDTH-1:0]   prod                ;
  logic signed  [WH_DATA_WIDTH-1:0]   prod_reg            ;

  logic         [ROW_LEN_WIDTH:0]     cnt                 ;

  logic                               calc_ena            ;
  logic                               calc_ena_reg        ;

  logic         [NUM_NODE_WIDTH-1:0]  num_node            ;
  logic         [NUM_NODE_WIDTH-1:0]  num_node_reg        ;
  logic         [NUM_NODE_WIDTH-1:0]  num_node_reg_q1     ;
  logic                               src_flag            ;
  logic                               src_flag_reg        ;
  logic                               src_flag_reg_q1     ;
  //* =========================================================

  integer i;

  //* =================== output assignment ===================
  assign res_o    = res_reg;
  assign pe_rdy_o = pe_rdy_reg;
  //* =========================================================


  //* ====================== calculation ======================
  assign wgt_addrb  = col_idx_i;
  assign calc_ena   = spmm_vld_q1;

  always_comb begin
    prod  = prod_reg;
    res   = res_reg;
    cnt   = cnt_reg;

    if (calc_ena_reg) begin
      prod  = wgt_dout;
      res   = (cnt_reg != 0) ? ($signed(res_reg) + $signed(wgt_dout)) : $signed(wgt_dout);
      cnt   = (cnt_reg == row_len_reg - 1 || row_len_reg <= 1) ? 0 : (cnt_reg + 1);
    end
  end

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      prod_reg      <= 'b0;
      cnt_reg       <= 'b0;
      res_reg       <= 'b0;
      calc_ena_reg  <= 'b0;
    end else begin
      cnt_reg       <= cnt;
      prod_reg      <= prod;
      res_reg       <= res;
      calc_ena_reg  <= calc_ena;
    end
  end

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      row_len_reg <= '0;
      spmm_vld_q1 <= '0;
    end else begin
      row_len_reg <= row_len_i;
      spmm_vld_q1 <= spmm_vld_i;
    end
  end
  //* =========================================================


  //* ======================== pe_rdy =========================
  always_comb begin
    pe_rdy = pe_rdy_reg;
    if (pe_rdy_reg && (row_len_reg > 1)) begin
      pe_rdy = 1'b0;
    end else if ((cnt_reg == row_len_reg - 1) || (row_len_reg == 1) && spmm_vld_i) begin
      pe_rdy = 1'b1;
    end
  end

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      pe_rdy_reg <= 'b0;
    end else begin
      if (row_len_reg == 1 && spmm_vld_i) begin
        pe_rdy_reg <= 1'b1;
      end else begin
        pe_rdy_reg <= pe_rdy;
      end
    end
  end
  //* =========================================================


  //* ======================= node_info =======================
  assign num_node_o = num_node_reg_q1;
  assign src_flag_o = src_flag_reg_q1;

  assign num_node = (pe_vld_i) ? num_node_i : num_node_reg;
  assign src_flag = (pe_vld_i) ? src_flag_i : src_flag_reg;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      num_node_reg    <= 'b0;
      num_node_reg_q1 <= 'b0;
      src_flag_reg    <= 'b0;
      src_flag_reg_q1 <= 'b0;
    end else begin
      num_node_reg    <= num_node;
      num_node_reg_q1 <= num_node_reg;
      src_flag_reg    <= src_flag;
      src_flag_reg_q1 <= src_flag_reg;
    end
  end
  //* =========================================================
endmodule