module aggregator #(

)(

);
endmodule